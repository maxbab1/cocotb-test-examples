// here it would be possible to instanciate multiple modules 
// to allow a testbench to test module interface compatibility
